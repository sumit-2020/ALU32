`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:34:56 12/07/2016 
// Design Name: 
// Module Name:    KoggeStone 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module KoggeStone(a,b,cin,sum,cout);
input [31:0] a,b;
input cin;
output [31:0] sum;
output cout;

	wire b1_2_gen, b1_2_prop;
	wire b1_3_gen, b1_3_prop;
	wire b1_4_gen, b1_4_prop;
	wire b1_5_gen, b1_5_prop;
	wire b1_6_gen, b1_6_prop;
	wire b1_7_gen, b1_7_prop;
	wire b1_8_gen, b1_8_prop;
	wire b1_9_gen, b1_9_prop;
	wire b1_10_gen, b1_10_prop;
	wire b1_11_gen, b1_11_prop;
	wire b1_12_gen, b1_12_prop;
	wire b1_13_gen, b1_13_prop;
	wire b1_14_gen, b1_14_prop;
	wire b1_15_gen, b1_15_prop;
	wire b1_16_gen, b1_16_prop;
	wire b1_17_gen, b1_17_prop;
	wire b1_18_gen, b1_18_prop;
	wire b1_19_gen, b1_19_prop;
	wire b1_20_gen, b1_20_prop;
	wire b1_21_gen, b1_21_prop;
	wire b1_22_gen, b1_22_prop;
	wire b1_23_gen, b1_23_prop;
	wire b1_24_gen, b1_24_prop;
	wire b1_25_gen, b1_25_prop;
	wire b1_26_gen, b1_26_prop;
	wire b1_27_gen, b1_27_prop;
	wire b1_28_gen, b1_28_prop;
	wire b1_29_gen, b1_29_prop;
	wire b1_30_gen, b1_30_prop;
	wire b1_31_gen, b1_31_prop;
	wire b2_4_gen, b2_4_prop;
	wire b2_5_gen, b2_5_prop;
	wire b2_6_gen, b2_6_prop;
	wire b2_7_gen, b2_7_prop;
	wire b2_8_gen, b2_8_prop;
	wire b2_9_gen, b2_9_prop;
	wire b2_10_gen, b2_10_prop;
	wire b2_11_gen, b2_11_prop;
	wire b2_12_gen, b2_12_prop;
	wire b2_13_gen, b2_13_prop;
	wire b2_14_gen, b2_14_prop;
	wire b2_15_gen, b2_15_prop;
	wire b2_16_gen, b2_16_prop;
	wire b2_17_gen, b2_17_prop;
	wire b2_18_gen, b2_18_prop;
	wire b2_19_gen, b2_19_prop;
	wire b2_20_gen, b2_20_prop;
	wire b2_21_gen, b2_21_prop;
	wire b2_22_gen, b2_22_prop;
	wire b2_23_gen, b2_23_prop;
	wire b2_24_gen, b2_24_prop;
	wire b2_25_gen, b2_25_prop;
	wire b2_26_gen, b2_26_prop;
	wire b2_27_gen, b2_27_prop;
	wire b2_28_gen, b2_28_prop;
	wire b2_29_gen, b2_29_prop;
	wire b2_30_gen, b2_30_prop;
	wire b2_31_gen, b2_31_prop;
	wire b3_8_gen, b3_8_prop;
	wire b3_9_gen, b3_9_prop;
	wire b3_10_gen, b3_10_prop;
	wire b3_11_gen, b3_11_prop;
	wire b3_12_gen, b3_12_prop;
	wire b3_13_gen, b3_13_prop;
	wire b3_14_gen, b3_14_prop;
	wire b3_15_gen, b3_15_prop;
	wire b3_16_gen, b3_16_prop;
	wire b3_17_gen, b3_17_prop;
	wire b3_18_gen, b3_18_prop;
	wire b3_19_gen, b3_19_prop;
	wire b3_20_gen, b3_20_prop;
	wire b3_21_gen, b3_21_prop;
	wire b3_22_gen, b3_22_prop;
	wire b3_23_gen, b3_23_prop;
	wire b3_24_gen, b3_24_prop;
	wire b3_25_gen, b3_25_prop;
	wire b3_26_gen, b3_26_prop;
	wire b3_27_gen, b3_27_prop;
	wire b3_28_gen, b3_28_prop;
	wire b3_29_gen, b3_29_prop;
	wire b3_30_gen, b3_30_prop;
	wire b3_31_gen, b3_31_prop;
	wire b4_16_gen, b4_16_prop;
	wire b4_17_gen, b4_17_prop;
	wire b4_18_gen, b4_18_prop;
	wire b4_19_gen, b4_19_prop;
	wire b4_20_gen, b4_20_prop;
	wire b4_21_gen, b4_21_prop;
	wire b4_22_gen, b4_22_prop;
	wire b4_23_gen, b4_23_prop;
	wire b4_24_gen, b4_24_prop;
	wire b4_25_gen, b4_25_prop;
	wire b4_26_gen, b4_26_prop;
	wire b4_27_gen, b4_27_prop;
	wire b4_28_gen, b4_28_prop;
	wire b4_29_gen, b4_29_prop;
	wire b4_30_gen, b4_30_prop;
	wire b4_31_gen, b4_31_prop;

wire g1_0_gen;
	assign g1_0_gen = cin;
	wire g1_1_gen;
	wire g2_2_gen;
	wire g2_3_gen;
	wire g3_4_gen;
	wire g3_5_gen;
	wire g3_6_gen;
	wire g3_7_gen;
	wire g4_8_gen;
	wire g4_9_gen;
	wire g4_10_gen;
	wire g4_11_gen;
	wire g4_12_gen;
	wire g4_13_gen;
	wire g4_14_gen;
	wire g4_15_gen;
	wire g5_16_gen;
	wire g5_17_gen;
	wire g5_18_gen;
	wire g5_19_gen;
	wire g5_20_gen;
	wire g5_21_gen;
	wire g5_22_gen;
	wire g5_23_gen;
	wire g5_24_gen;
	wire g5_25_gen;
	wire g5_26_gen;
	wire g5_27_gen;
	wire g5_28_gen;
	wire g5_29_gen;
	wire g5_30_gen;
	wire g5_31_gen;
	
	wire [31:0] gen,prop;

	assign gen[0]=cin;
	assign prop[0]=1'b1;
	GP gp1(a[0], b[0] , gen[1], prop[1]);
	GP gp2(a[1], b[1] , gen[2], prop[2]);
	GP gp3(a[2], b[2] , gen[3], prop[3]);
	GP gp4(a[3], b[3] , gen[4], prop[4]);
	GP gp5(a[4], b[4] , gen[5], prop[5]);
	GP gp6(a[5], b[5] , gen[6], prop[6]);
	GP gp7(a[6], b[6] , gen[7], prop[7]);
	GP gp8(a[7], b[7] , gen[8], prop[8]);
	GP gp9(a[8], b[8] , gen[9], prop[9]);
	GP gp10(a[9], b[9] , gen[10], prop[10]);
	GP gp11(a[10], b[10] , gen[11], prop[11]);
	GP gp12(a[11], b[11] , gen[12], prop[12]);
	GP gp13(a[12], b[12] , gen[13], prop[13]);
	GP gp14(a[13], b[13] , gen[14], prop[14]);
	GP gp15(a[14], b[14] , gen[15], prop[15]);
	GP gp16(a[15], b[15] , gen[16], prop[16]);
	GP gp17(a[16], b[16] , gen[17], prop[17]);
	GP gp18(a[17], b[17] , gen[18], prop[18]);
	GP gp19(a[18], b[18] , gen[19], prop[19]);
	GP gp20(a[19], b[19] , gen[20], prop[20]);
	GP gp21(a[20], b[20] , gen[21], prop[21]);
	GP gp22(a[21], b[21] , gen[22], prop[22]);
	GP gp23(a[22], b[22] , gen[23], prop[23]);
	GP gp24(a[23], b[23] , gen[24], prop[24]);
	GP gp25(a[24], b[24] , gen[25], prop[25]);
	GP gp26(a[25], b[25] , gen[26], prop[26]);
	GP gp27(a[26], b[26] , gen[27], prop[27]);
	GP gp28(a[27], b[27] , gen[28], prop[28]);
	GP gp29(a[28], b[28] , gen[29], prop[29]);
	GP gp30(a[29], b[29] , gen[30], prop[30]);
	GP gp31(a[30], b[30] , gen[31], prop[31]);

	Black b1_2(gen[2], prop[2] , gen[1], prop[1], b1_2_gen, b1_2_prop);
	Black b1_3(gen[3], prop[3] , gen[2], prop[2], b1_3_gen, b1_3_prop);
	Black b1_4(gen[4], prop[4] , gen[3], prop[3], b1_4_gen, b1_4_prop);
	Black b1_5(gen[5], prop[5] , gen[4], prop[4], b1_5_gen, b1_5_prop);
	Black b1_6(gen[6], prop[6] , gen[5], prop[5], b1_6_gen, b1_6_prop);
	Black b1_7(gen[7], prop[7] , gen[6], prop[6], b1_7_gen, b1_7_prop);
	Black b1_8(gen[8], prop[8] , gen[7], prop[7], b1_8_gen, b1_8_prop);
	Black b1_9(gen[9], prop[9] , gen[8], prop[8], b1_9_gen, b1_9_prop);
	Black b1_10(gen[10], prop[10] , gen[9], prop[9], b1_10_gen, b1_10_prop);
	Black b1_11(gen[11], prop[11] , gen[10], prop[10], b1_11_gen, b1_11_prop);
	Black b1_12(gen[12], prop[12] , gen[11], prop[11], b1_12_gen, b1_12_prop);
	Black b1_13(gen[13], prop[13] , gen[12], prop[12], b1_13_gen, b1_13_prop);
	Black b1_14(gen[14], prop[14] , gen[13], prop[13], b1_14_gen, b1_14_prop);
	Black b1_15(gen[15], prop[15] , gen[14], prop[14], b1_15_gen, b1_15_prop);
	Black b1_16(gen[16], prop[16] , gen[15], prop[15], b1_16_gen, b1_16_prop);
	Black b1_17(gen[17], prop[17] , gen[16], prop[16], b1_17_gen, b1_17_prop);
	Black b1_18(gen[18], prop[18] , gen[17], prop[17], b1_18_gen, b1_18_prop);
	Black b1_19(gen[19], prop[19] , gen[18], prop[18], b1_19_gen, b1_19_prop);
	Black b1_20(gen[20], prop[20] , gen[19], prop[19], b1_20_gen, b1_20_prop);
	Black b1_21(gen[21], prop[21] , gen[20], prop[20], b1_21_gen, b1_21_prop);
	Black b1_22(gen[22], prop[22] , gen[21], prop[21], b1_22_gen, b1_22_prop);
	Black b1_23(gen[23], prop[23] , gen[22], prop[22], b1_23_gen, b1_23_prop);
	Black b1_24(gen[24], prop[24] , gen[23], prop[23], b1_24_gen, b1_24_prop);
	Black b1_25(gen[25], prop[25] , gen[24], prop[24], b1_25_gen, b1_25_prop);
	Black b1_26(gen[26], prop[26] , gen[25], prop[25], b1_26_gen, b1_26_prop);
	Black b1_27(gen[27], prop[27] , gen[26], prop[26], b1_27_gen, b1_27_prop);
	Black b1_28(gen[28], prop[28] , gen[27], prop[27], b1_28_gen, b1_28_prop);
	Black b1_29(gen[29], prop[29] , gen[28], prop[28], b1_29_gen, b1_29_prop);
	Black b1_30(gen[30], prop[30] , gen[29], prop[29], b1_30_gen, b1_30_prop);
	Black b1_31(gen[31], prop[31] , gen[30], prop[30], b1_31_gen, b1_31_prop);

	Black b2_4(b1_4_gen, b1_4_prop, b1_2_gen, b1_2_prop, b2_4_gen, b2_4_prop);
	Black b2_5(b1_5_gen, b1_5_prop, b1_3_gen, b1_3_prop, b2_5_gen, b2_5_prop);
	Black b2_6(b1_6_gen, b1_6_prop, b1_4_gen, b1_4_prop, b2_6_gen, b2_6_prop);
	Black b2_7(b1_7_gen, b1_7_prop, b1_5_gen, b1_5_prop, b2_7_gen, b2_7_prop);
	Black b2_8(b1_8_gen, b1_8_prop, b1_6_gen, b1_6_prop, b2_8_gen, b2_8_prop);
	Black b2_9(b1_9_gen, b1_9_prop, b1_7_gen, b1_7_prop, b2_9_gen, b2_9_prop);
	Black b2_10(b1_10_gen, b1_10_prop, b1_8_gen, b1_8_prop, b2_10_gen, b2_10_prop);
	Black b2_11(b1_11_gen, b1_11_prop, b1_9_gen, b1_9_prop, b2_11_gen, b2_11_prop);
	Black b2_12(b1_12_gen, b1_12_prop, b1_10_gen, b1_10_prop, b2_12_gen, b2_12_prop);
	Black b2_13(b1_13_gen, b1_13_prop, b1_11_gen, b1_11_prop, b2_13_gen, b2_13_prop);
	Black b2_14(b1_14_gen, b1_14_prop, b1_12_gen, b1_12_prop, b2_14_gen, b2_14_prop);
	Black b2_15(b1_15_gen, b1_15_prop, b1_13_gen, b1_13_prop, b2_15_gen, b2_15_prop);
	Black b2_16(b1_16_gen, b1_16_prop, b1_14_gen, b1_14_prop, b2_16_gen, b2_16_prop);
	Black b2_17(b1_17_gen, b1_17_prop, b1_15_gen, b1_15_prop, b2_17_gen, b2_17_prop);
	Black b2_18(b1_18_gen, b1_18_prop, b1_16_gen, b1_16_prop, b2_18_gen, b2_18_prop);
	Black b2_19(b1_19_gen, b1_19_prop, b1_17_gen, b1_17_prop, b2_19_gen, b2_19_prop);
	Black b2_20(b1_20_gen, b1_20_prop, b1_18_gen, b1_18_prop, b2_20_gen, b2_20_prop);
	Black b2_21(b1_21_gen, b1_21_prop, b1_19_gen, b1_19_prop, b2_21_gen, b2_21_prop);
	Black b2_22(b1_22_gen, b1_22_prop, b1_20_gen, b1_20_prop, b2_22_gen, b2_22_prop);
	Black b2_23(b1_23_gen, b1_23_prop, b1_21_gen, b1_21_prop, b2_23_gen, b2_23_prop);
	Black b2_24(b1_24_gen, b1_24_prop, b1_22_gen, b1_22_prop, b2_24_gen, b2_24_prop);
	Black b2_25(b1_25_gen, b1_25_prop, b1_23_gen, b1_23_prop, b2_25_gen, b2_25_prop);
	Black b2_26(b1_26_gen, b1_26_prop, b1_24_gen, b1_24_prop, b2_26_gen, b2_26_prop);
	Black b2_27(b1_27_gen, b1_27_prop, b1_25_gen, b1_25_prop, b2_27_gen, b2_27_prop);
	Black b2_28(b1_28_gen, b1_28_prop, b1_26_gen, b1_26_prop, b2_28_gen, b2_28_prop);
	Black b2_29(b1_29_gen, b1_29_prop, b1_27_gen, b1_27_prop, b2_29_gen, b2_29_prop);
	Black b2_30(b1_30_gen, b1_30_prop, b1_28_gen, b1_28_prop, b2_30_gen, b2_30_prop);
	Black b2_31(b1_31_gen, b1_31_prop, b1_29_gen, b1_29_prop, b2_31_gen, b2_31_prop);
	Black b3_8(b2_8_gen, b2_8_prop, b2_4_gen, b2_4_prop, b3_8_gen, b3_8_prop);
	Black b3_9(b2_9_gen, b2_9_prop, b2_5_gen, b2_5_prop, b3_9_gen, b3_9_prop);
	Black b3_10(b2_10_gen, b2_10_prop, b2_6_gen, b2_6_prop, b3_10_gen, b3_10_prop);
	Black b3_11(b2_11_gen, b2_11_prop, b2_7_gen, b2_7_prop, b3_11_gen, b3_11_prop);
	Black b3_12(b2_12_gen, b2_12_prop, b2_8_gen, b2_8_prop, b3_12_gen, b3_12_prop);
	Black b3_13(b2_13_gen, b2_13_prop, b2_9_gen, b2_9_prop, b3_13_gen, b3_13_prop);
	Black b3_14(b2_14_gen, b2_14_prop, b2_10_gen, b2_10_prop, b3_14_gen, b3_14_prop);
	Black b3_15(b2_15_gen, b2_15_prop, b2_11_gen, b2_11_prop, b3_15_gen, b3_15_prop);
	Black b3_16(b2_16_gen, b2_16_prop, b2_12_gen, b2_12_prop, b3_16_gen, b3_16_prop);
	Black b3_17(b2_17_gen, b2_17_prop, b2_13_gen, b2_13_prop, b3_17_gen, b3_17_prop);
	Black b3_18(b2_18_gen, b2_18_prop, b2_14_gen, b2_14_prop, b3_18_gen, b3_18_prop);
	Black b3_19(b2_19_gen, b2_19_prop, b2_15_gen, b2_15_prop, b3_19_gen, b3_19_prop);
	Black b3_20(b2_20_gen, b2_20_prop, b2_16_gen, b2_16_prop, b3_20_gen, b3_20_prop);
	Black b3_21(b2_21_gen, b2_21_prop, b2_17_gen, b2_17_prop, b3_21_gen, b3_21_prop);
	Black b3_22(b2_22_gen, b2_22_prop, b2_18_gen, b2_18_prop, b3_22_gen, b3_22_prop);
	Black b3_23(b2_23_gen, b2_23_prop, b2_19_gen, b2_19_prop, b3_23_gen, b3_23_prop);
	Black b3_24(b2_24_gen, b2_24_prop, b2_20_gen, b2_20_prop, b3_24_gen, b3_24_prop);
	Black b3_25(b2_25_gen, b2_25_prop, b2_21_gen, b2_21_prop, b3_25_gen, b3_25_prop);
	Black b3_26(b2_26_gen, b2_26_prop, b2_22_gen, b2_22_prop, b3_26_gen, b3_26_prop);
	Black b3_27(b2_27_gen, b2_27_prop, b2_23_gen, b2_23_prop, b3_27_gen, b3_27_prop);
	Black b3_28(b2_28_gen, b2_28_prop, b2_24_gen, b2_24_prop, b3_28_gen, b3_28_prop);
	Black b3_29(b2_29_gen, b2_29_prop, b2_25_gen, b2_25_prop, b3_29_gen, b3_29_prop);
	Black b3_30(b2_30_gen, b2_30_prop, b2_26_gen, b2_26_prop, b3_30_gen, b3_30_prop);
	Black b3_31(b2_31_gen, b2_31_prop, b2_27_gen, b2_27_prop, b3_31_gen, b3_31_prop);
	Black b4_16(b3_16_gen, b3_16_prop, b3_8_gen, b3_8_prop, b4_16_gen, b4_16_prop);
	Black b4_17(b3_17_gen, b3_17_prop, b3_9_gen, b3_9_prop, b4_17_gen, b4_17_prop);
	Black b4_18(b3_18_gen, b3_18_prop, b3_10_gen, b3_10_prop, b4_18_gen, b4_18_prop);
	Black b4_19(b3_19_gen, b3_19_prop, b3_11_gen, b3_11_prop, b4_19_gen, b4_19_prop);
	Black b4_20(b3_20_gen, b3_20_prop, b3_12_gen, b3_12_prop, b4_20_gen, b4_20_prop);
	Black b4_21(b3_21_gen, b3_21_prop, b3_13_gen, b3_13_prop, b4_21_gen, b4_21_prop);
	Black b4_22(b3_22_gen, b3_22_prop, b3_14_gen, b3_14_prop, b4_22_gen, b4_22_prop);
	Black b4_23(b3_23_gen, b3_23_prop, b3_15_gen, b3_15_prop, b4_23_gen, b4_23_prop);
	Black b4_24(b3_24_gen, b3_24_prop, b3_16_gen, b3_16_prop, b4_24_gen, b4_24_prop);
	Black b4_25(b3_25_gen, b3_25_prop, b3_17_gen, b3_17_prop, b4_25_gen, b4_25_prop);
	Black b4_26(b3_26_gen, b3_26_prop, b3_18_gen, b3_18_prop, b4_26_gen, b4_26_prop);
	Black b4_27(b3_27_gen, b3_27_prop, b3_19_gen, b3_19_prop, b4_27_gen, b4_27_prop);
	Black b4_28(b3_28_gen, b3_28_prop, b3_20_gen, b3_20_prop, b4_28_gen, b4_28_prop);
	Black b4_29(b3_29_gen, b3_29_prop, b3_21_gen, b3_21_prop, b4_29_gen, b4_29_prop);
	Black b4_30(b3_30_gen, b3_30_prop, b3_22_gen, b3_22_prop, b4_30_gen, b4_30_prop);
	Black b4_31(b3_31_gen, b3_31_prop, b3_23_gen, b3_23_prop, b4_31_gen, b4_31_prop);

	Grey g1_1(gen[1], prop[1], cin, g1_1_gen);
	Grey g2_2(b1_2_gen, b1_2_prop, cin, g2_2_gen);
	Grey g2_3(b1_3_gen, b1_3_prop, g1_1_gen, g2_3_gen);
	Grey g3_4(b2_4_gen, b2_4_prop, cin, g3_4_gen);
	Grey g3_5(b2_5_gen, b2_5_prop, g1_1_gen, g3_5_gen);
	Grey g3_6(b2_6_gen, b2_6_prop, g2_2_gen, g3_6_gen);
	Grey g3_7(b2_7_gen, b2_7_prop, g2_3_gen, g3_7_gen);
	Grey g4_8(b3_8_gen, b3_8_prop, cin, g4_8_gen);
	Grey g4_9(b3_9_gen, b3_9_prop, g1_1_gen, g4_9_gen);
	Grey g4_10(b3_10_gen, b3_10_prop, g2_2_gen, g4_10_gen);
	Grey g4_11(b3_11_gen, b3_11_prop, g2_3_gen, g4_11_gen);
	Grey g4_12(b3_12_gen, b3_12_prop, g3_4_gen, g4_12_gen);
	Grey g4_13(b3_13_gen, b3_13_prop, g3_5_gen, g4_13_gen);
	Grey g4_14(b3_14_gen, b3_14_prop, g3_6_gen, g4_14_gen);
	Grey g4_15(b3_15_gen, b3_15_prop, g3_7_gen, g4_15_gen);
	Grey g5_16(b4_16_gen, b4_16_prop, cin, g5_16_gen);
	Grey g5_17(b4_17_gen, b4_17_prop, g1_1_gen, g5_17_gen);
	Grey g5_18(b4_18_gen, b4_18_prop, g2_2_gen, g5_18_gen);
	Grey g5_19(b4_19_gen, b4_19_prop, g2_3_gen, g5_19_gen);
	Grey g5_20(b4_20_gen, b4_20_prop, g3_4_gen, g5_20_gen);
	Grey g5_21(b4_21_gen, b4_21_prop, g3_5_gen, g5_21_gen);
	Grey g5_22(b4_22_gen, b4_22_prop, g3_6_gen, g5_22_gen);
	Grey g5_23(b4_23_gen, b4_23_prop, g3_7_gen, g5_23_gen);
	Grey g5_24(b4_24_gen, b4_24_prop, g4_8_gen, g5_24_gen);
	Grey g5_25(b4_25_gen, b4_25_prop, g4_9_gen, g5_25_gen);
	Grey g5_26(b4_26_gen, b4_26_prop, g4_10_gen, g5_26_gen);
	Grey g5_27(b4_27_gen, b4_27_prop, g4_11_gen, g5_27_gen);
	Grey g5_28(b4_28_gen, b4_28_prop, g4_12_gen, g5_28_gen);
	Grey g5_29(b4_29_gen, b4_29_prop, g4_13_gen, g5_29_gen);
	Grey g5_30(b4_30_gen, b4_30_prop, g4_14_gen, g5_30_gen);
	Grey g5_31(b4_31_gen, b4_31_prop, g4_15_gen, g5_31_gen);
	
	xor(sum[0],a[0]^b[0],cin);
	xor(sum[1], prop[2], g1_1_gen);
	xor(sum[2], prop[3], g2_2_gen);
	xor(sum[3], prop[4], g2_3_gen);
	xor(sum[4], prop[5], g3_4_gen);
	xor(sum[5], prop[6], g3_5_gen);
	xor(sum[6], prop[7], g3_6_gen);
	xor(sum[7], prop[8], g3_7_gen);
	xor(sum[8], prop[9], g4_8_gen);
	xor(sum[9], prop[10], g4_9_gen);
	xor(sum[10], prop[11], g4_10_gen);
	xor(sum[11], prop[12], g4_11_gen);
	xor(sum[12], prop[13], g4_12_gen);
	xor(sum[13], prop[14], g4_13_gen);
	xor(sum[14], prop[15], g4_14_gen);
	xor(sum[15], prop[16], g4_15_gen);
	xor(sum[16], prop[17], g5_16_gen);
	xor(sum[17], prop[18], g5_17_gen);
	xor(sum[18], prop[19], g5_18_gen);
	xor(sum[19], prop[20], g5_19_gen);
	xor(sum[20], prop[21], g5_20_gen);
	xor(sum[21], prop[22], g5_21_gen);
	xor(sum[22], prop[23], g5_22_gen);
	xor(sum[23], prop[24], g5_23_gen);
	xor(sum[24], prop[25], g5_24_gen);
	xor(sum[25], prop[26], g5_25_gen);
	xor(sum[26], prop[27], g5_26_gen);
	xor(sum[27], prop[28], g5_27_gen);
	xor(sum[28], prop[29], g5_28_gen);
	xor(sum[29], prop[30], g5_29_gen);
	xor(sum[30], prop[31], g5_30_gen);
	xor(sum[31], a[31]^b[31], g5_31_gen);

	wire temp=prop[31]*g5_31_gen;
	or(cout,gen[31],temp);


endmodule
